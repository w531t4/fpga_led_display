`default_nettype none
(* blackbox *)
module EHXPLLL (
        input CLKI, CLKFB,
        input PHASESEL1, PHASESEL0, PHASEDIR, PHASESTEP, PHASELOADREG,
        input STDBY, PLLWAKESYNC,
        input RST, ENCLKOP, ENCLKOS, ENCLKOS2, ENCLKOS3,
        output CLKOP, CLKOS, CLKOS2, CLKOS3,
        output LOCK, INTLOCK,
        output REFCLK, CLKINTFB
);
        parameter CLKI_DIV = 1;
        parameter CLKFB_DIV = 1;
        parameter CLKOP_DIV = 8;
        parameter CLKOS_DIV = 8;
        parameter CLKOS2_DIV = 8;
        parameter CLKOS3_DIV = 8;
        parameter CLKOP_ENABLE = "ENABLED";
        parameter CLKOS_ENABLE = "DISABLED";
        parameter CLKOS2_ENABLE = "DISABLED";
        parameter CLKOS3_ENABLE = "DISABLED";
        parameter CLKOP_CPHASE = 0;
        parameter CLKOS_CPHASE = 0;
        parameter CLKOS2_CPHASE = 0;
        parameter CLKOS3_CPHASE = 0;
        parameter CLKOP_FPHASE = 0;
        parameter CLKOS_FPHASE = 0;
        parameter CLKOS2_FPHASE = 0;
        parameter CLKOS3_FPHASE = 0;
        parameter FEEDBK_PATH = "CLKOP";
        parameter CLKOP_TRIM_POL = "RISING";
        parameter CLKOP_TRIM_DELAY = 0;
        parameter CLKOS_TRIM_POL = "RISING";
        parameter CLKOS_TRIM_DELAY = 0;
        parameter OUTDIVIDER_MUXA = "DIVA";
        parameter OUTDIVIDER_MUXB = "DIVB";
        parameter OUTDIVIDER_MUXC = "DIVC";
        parameter OUTDIVIDER_MUXD = "DIVD";
        parameter PLL_LOCK_MODE = 0;
        parameter PLL_LOCK_DELAY = 200;
        parameter STDBY_ENABLE = "DISABLED";
        parameter REFIN_RESET = "DISABLED";
        parameter SYNC_ENABLE = "DISABLED";
        parameter INT_LOCK_STICKY = "ENABLED";
        parameter DPHASE_SOURCE = "DISABLED";
        parameter PLLRST_ENA = "DISABLED";
        parameter INTFB_WAKE = "DISABLED";
endmodule

module DP16KD(
  input DIA17, DIA16, DIA15, DIA14, DIA13, DIA12, DIA11, DIA10, DIA9, DIA8, DIA7, DIA6, DIA5, DIA4, DIA3, DIA2, DIA1, DIA0,
  input ADA13, ADA12, ADA11, ADA10, ADA9, ADA8, ADA7, ADA6, ADA5, ADA4, ADA3, ADA2, ADA1, ADA0,
  input CEA, OCEA, CLKA, WEA, RSTA,
  input CSA2, CSA1, CSA0,
  output DOA17, DOA16, DOA15, DOA14, DOA13, DOA12, DOA11, DOA10, DOA9, DOA8, DOA7, DOA6, DOA5, DOA4, DOA3, DOA2, DOA1, DOA0,

  input DIB17, DIB16, DIB15, DIB14, DIB13, DIB12, DIB11, DIB10, DIB9, DIB8, DIB7, DIB6, DIB5, DIB4, DIB3, DIB2, DIB1, DIB0,
  input ADB13, ADB12, ADB11, ADB10, ADB9, ADB8, ADB7, ADB6, ADB5, ADB4, ADB3, ADB2, ADB1, ADB0,
  input CEB, OCEB, CLKB, WEB, RSTB,
  input CSB2, CSB1, CSB0,
  output DOB17, DOB16, DOB15, DOB14, DOB13, DOB12, DOB11, DOB10, DOB9, DOB8, DOB7, DOB6, DOB5, DOB4, DOB3, DOB2, DOB1, DOB0
);
        parameter DATA_WIDTH_A = 18;
        parameter DATA_WIDTH_B = 18;

        parameter REGMODE_A = "NOREG";
        parameter REGMODE_B = "NOREG";

        parameter RESETMODE = "SYNC";
        parameter ASYNC_RESET_RELEASE = "SYNC";

        parameter CSDECODE_A = "0b000";
        parameter CSDECODE_B = "0b000";

        parameter WRITEMODE_A = "NORMAL";
        parameter WRITEMODE_B = "NORMAL";

        parameter DIA17MUX = "DIA17";
        parameter DIA16MUX = "DIA16";
        parameter DIA15MUX = "DIA15";
        parameter DIA14MUX = "DIA14";
        parameter DIA13MUX = "DIA13";
        parameter DIA12MUX = "DIA12";
        parameter DIA11MUX = "DIA11";
        parameter DIA10MUX = "DIA10";
        parameter DIA9MUX = "DIA9";
        parameter DIA8MUX = "DIA8";
        parameter DIA7MUX = "DIA7";
        parameter DIA6MUX = "DIA6";
        parameter DIA5MUX = "DIA5";
        parameter DIA4MUX = "DIA4";
        parameter DIA3MUX = "DIA3";
        parameter DIA2MUX = "DIA2";
        parameter DIA1MUX = "DIA1";
        parameter DIA0MUX = "DIA0";
        parameter ADA13MUX = "ADA13";
        parameter ADA12MUX = "ADA12";
        parameter ADA11MUX = "ADA11";
        parameter ADA10MUX = "ADA10";
        parameter ADA9MUX = "ADA9";
        parameter ADA8MUX = "ADA8";
        parameter ADA7MUX = "ADA7";
        parameter ADA6MUX = "ADA6";
        parameter ADA5MUX = "ADA5";
        parameter ADA4MUX = "ADA4";
        parameter ADA3MUX = "ADA3";
        parameter ADA2MUX = "ADA2";
        parameter ADA1MUX = "ADA1";
        parameter ADA0MUX = "ADA0";
        parameter CEAMUX = "CEA";
        parameter OCEAMUX = "OCEA";
        parameter CLKAMUX = "CLKA";
        parameter WEAMUX = "WEA";
        parameter RSTAMUX = "RSTA";
        parameter CSA2MUX = "CSA2";
        parameter CSA1MUX = "CSA1";
        parameter CSA0MUX = "CSA0";
        parameter DOA17MUX = "DOA17";
        parameter DOA16MUX = "DOA16";
        parameter DOA15MUX = "DOA15";
        parameter DOA14MUX = "DOA14";
        parameter DOA13MUX = "DOA13";
        parameter DOA12MUX = "DOA12";
        parameter DOA11MUX = "DOA11";
        parameter DOA10MUX = "DOA10";
        parameter DOA9MUX = "DOA9";
        parameter DOA8MUX = "DOA8";
        parameter DOA7MUX = "DOA7";
        parameter DOA6MUX = "DOA6";
        parameter DOA5MUX = "DOA5";
        parameter DOA4MUX = "DOA4";
        parameter DOA3MUX = "DOA3";
        parameter DOA2MUX = "DOA2";
        parameter DOA1MUX = "DOA1";
        parameter DOA0MUX = "DOA0";
        parameter DIB17MUX = "DIB17";
        parameter DIB16MUX = "DIB16";
        parameter DIB15MUX = "DIB15";
        parameter DIB14MUX = "DIB14";
        parameter DIB13MUX = "DIB13";
        parameter DIB12MUX = "DIB12";
        parameter DIB11MUX = "DIB11";
        parameter DIB10MUX = "DIB10";
        parameter DIB9MUX = "DIB9";
        parameter DIB8MUX = "DIB8";
        parameter DIB7MUX = "DIB7";
        parameter DIB6MUX = "DIB6";
        parameter DIB5MUX = "DIB5";
        parameter DIB4MUX = "DIB4";
        parameter DIB3MUX = "DIB3";
        parameter DIB2MUX = "DIB2";
        parameter DIB1MUX = "DIB1";
        parameter DIB0MUX = "DIB0";
        parameter ADB13MUX = "ADB13";
        parameter ADB12MUX = "ADB12";
        parameter ADB11MUX = "ADB11";
        parameter ADB10MUX = "ADB10";
        parameter ADB9MUX = "ADB9";
        parameter ADB8MUX = "ADB8";
        parameter ADB7MUX = "ADB7";
        parameter ADB6MUX = "ADB6";
        parameter ADB5MUX = "ADB5";
        parameter ADB4MUX = "ADB4";
        parameter ADB3MUX = "ADB3";
        parameter ADB2MUX = "ADB2";
        parameter ADB1MUX = "ADB1";
        parameter ADB0MUX = "ADB0";
        parameter CEBMUX = "CEB";
        parameter OCEBMUX = "OCEB";
        parameter CLKBMUX = "CLKB";
        parameter WEBMUX = "WEB";
        parameter RSTBMUX = "RSTB";
        parameter CSB2MUX = "CSB2";
        parameter CSB1MUX = "CSB1";
        parameter CSB0MUX = "CSB0";
        parameter DOB17MUX = "DOB17";
        parameter DOB16MUX = "DOB16";
        parameter DOB15MUX = "DOB15";
        parameter DOB14MUX = "DOB14";
        parameter DOB13MUX = "DOB13";
        parameter DOB12MUX = "DOB12";
        parameter DOB11MUX = "DOB11";
        parameter DOB10MUX = "DOB10";
        parameter DOB9MUX = "DOB9";
        parameter DOB8MUX = "DOB8";
        parameter DOB7MUX = "DOB7";
        parameter DOB6MUX = "DOB6";
        parameter DOB5MUX = "DOB5";
        parameter DOB4MUX = "DOB4";
        parameter DOB3MUX = "DOB3";
        parameter DOB2MUX = "DOB2";
        parameter DOB1MUX = "DOB1";
        parameter DOB0MUX = "DOB0";

        parameter WID = 0;

        parameter GSR = "ENABLED";

        parameter INITVAL_00 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_01 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_02 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_03 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_04 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_05 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_06 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_07 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_08 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_09 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_0A = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_0B = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_0C = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_0D = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_0E = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_0F = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_10 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_11 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_12 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_13 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_14 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_15 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_16 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_17 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_18 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_19 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_1A = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_1B = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_1C = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_1D = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_1E = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_1F = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_20 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_21 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_22 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_23 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_24 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_25 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_26 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_27 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_28 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_29 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_2A = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_2B = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_2C = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_2D = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_2E = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_2F = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_30 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_31 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_32 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_33 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_34 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_35 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_36 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_37 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_38 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_39 = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_3A = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_3B = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_3C = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_3D = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_3E = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INITVAL_3F = 320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000;
        parameter INIT_DATA = "STATIC";
endmodule

module VLO(output Z);
        assign Z = 1'b0;
endmodule

module VHI(output Z);
        assign Z = 1'b1;
endmodule

(* blackbox, keep *)
module GSR (
        input GSR
);
endmodule

(* blackbox *)
module PUR (
        input PUR
);
        parameter RST_PULSE = 1;
endmodule


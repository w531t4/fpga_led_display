`ifdef JUNK
    //>>> "".join([a[i] for i in range(len(a)-1, -1, -1)])
    //'brR L-77665544332211887766554433221188776655443322118877665544332211887766554433221188776655443322118877665544332211887766554433221110'
    //logic [1071:0] mystring = "brR L-77665544332211887766554433221188776655443322118877665544332211887766554433221188776655443322118877665544332211887766554433221110";
    //logic [1071:0] mystring = 'h627252204c2d3737363635353434333332323131383837373636353534343333323231313838373736363535343433333232313138383737363635353434333332323131383837373636353534343333323231313838373736363535343433333232313138383737363635353434333332323131383837373636353534343333323231313130;
    //logic [2111:0] mystring = 'h627252204c2d37373636353534343333323231313838373736363535343433333232313138383737363635353434333332323131383837373636353534343333323231313838373736363535343433333232313138383737363635353434333332323131383837373636353534343333323231313838373736363535343433333232313131304c133737363635353434333332323131383837373636353534343333323231313838373736363535343433333232313138383737363635353434333332323131383837373636353534343333323231313838373736363535343433333232313138383737363635353434333332323131383837373636353534343333323231313130;

    // switched 4c18 to 4c09 (in an effort to align 4c09 with 4c19 [which immediately follows])
    // for some reason this seems to start simulating at 4c18 (row 22..)
    // also, for 4c09 added 0x1234 as first few pixels, and for 4c19 added 0x5678 for first few pixels
    // 8320 * 8 = 66560, log2=16.001... -> 17
    // mystring represents many concatenated led pixel rows (L01DATA,L02DATA...)
    // logic [66559:0] mystringfull = 'h4c0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004c0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004c0200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004c030000000000009800980098000000000081a081a081a081a000000000000094c094c094c000000000042004200420042000000000044f044f044f044f044f0000021002100210021002100000000000160016001600000000401300000000000040130000881188118811881188110000000000009800980098000000000000004c040000000098000000000000009800000081a000000000000081a0000094c000000000000094c00000042000000000000004200000044f00000000000000000000021000000000000000000000001600000000000000160000401300000000000040130000000000008811000000000000000000000000980000000000000000004c050000000098000000000000009800000081a000000000000081a0000094c000000000000000000000042000000000000004200000044f00000000000000000000021000000000000000000000001600000000000000000000401300000000000040130000000000008811000000000000000000000000980000000000000000004c060000000098000000000000009800000081a081a081a081a00000000094c000000000000000000000042000000000000004200000044f044f044f044f00000000021002100210021000000000001600000000000000000000401340134013401340130000000000008811000000000000000000000000980000000000000000004c070000000098009800980098009800000081a000000000000081a0000094c000000000000000000000042000000000000004200000044f00000000000000000000021000000000000000000000001600000000001600160000401300000000000040130000000000008811000000000000000000000000980000000000000000004c080000000098000000000000009800000081a000000000000081a0000094c000000000000094c00000042000000000000004200000044f00000000000000000000021000000000000000000000001600000000000000160000401300000000000040130000000000008811000000000000980000000000980000000000000000004c090000000098000000000000009800000081a081a081a081a000000000000094c094c094c000000000042004200420042000000000044f044f044f044f044f0000021000000000000000000000000000160016001600000000401300000000000040130000881188118811881188110000000098009800000000000000000000004c0a00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004c0b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004c0c00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004c0d00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004c0e0000000000000000000000000000000081a000000000000000000000000000000000000000000000000000000000000004200000000000000000000000000000000000000210021000000000000000000000000000000000401300000000000000000000000000008811000000000000000000000000980000000000000000004c0f0000000000000000000000000000000081a000000000000000000000000000000000000000000000000000000000000004200000000000000000000000000000000002100000000002100000000000000000000000000000401300000000000000000000000000000000000000000000000000000000000000000000000000004c100000000000009800980098000000000081a0000081a081a000000000000094c094c094c0000000000000042004200000042000000000044f044f044f00000000000002100000000000000000000000160016001600160000401300004013401300000000000000008811000000000000000000009800980000000000000000004c110000000000000000000000009800000081a081a00000000081a0000094c000000000000000000000042000000000042004200000044f000000000000044f0000021002100210000000000000001600000000000000160000401340130000000040130000000088118811000000000000000000000000980000000000000000004c120000000000009800980098009800000081a000000000000081a0000094c000000000000000000000042000000000000004200000044f044f044f044f00000000000002100000000000000000000000160016001600160000401300000000000040130000000000008811000000000000000000000000980000000000000000004c130000000098000000000000009800000081a000000000000081a0000094c000000000000094c00000042000000000000004200000044f00000000000000000000000002100000000000000000000000000000000000160000401300000000000040130000000000008811000000000000980000000000980000000000000000004c140000000000009800980098000000000081a081a081a081a000000000000094c094c094c0000000000000042004200420042000000000044f044f044f00000000000002100000000000000000000000160016001600000000401300000000000040130000000088118811881100000000000098009800000000000000000000004c1500000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004c1600000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004c17000000000000980098009800000000000000000081a0000000000000000094c094c094c000000000042004200420042004200000000000000000044f00000000021002100210021002100000000000000016001600000000401340134013401340130000000088118811881100000000000098009800980000000000000000004c0912340000980000000000000098000000000081a081a000000000000094c000000000000094c0000000000000000004200000000000000000044f044f00000000021000000000000000000000000000160000000000000000401300000000000040130000881100000000000088110000980000000000000098000000000000004c19567800009800000000009800980000000000000081a0000000000000000000000000000094c00000000000000420000000000000000002100000044f00000000021002100210021000000000001600000000000000000000000000000000401300000000881100000000000088110000980000000000000098000000000000004c1a000000009800000098000000980000000000000081a000000000000000000000000094c000000000000000000000042000000000044f00000000044f00000000000000000000000002100000001600160016001600000000000000000000401300000000000088118811881100000000000098009800980098000000000000004c1b000000009800980000000000980000000000000081a00000000000000000000094c0000000000000000000000000000004200000044f044f044f044f044f0000000000000000000002100000001600000000000000160000000000004013000000000000881100000000000088110000000000000000000098000000000000004c1c000000009800000000000000980000000000000081a0000000000000000094c00000000000000000042000000000000004200000000000000000044f00000000021000000000000002100000001600000000000000160000000000004013000000000000881100000000000088110000000000000000980000000000000000004c1d00000000000098009800980000000000000081a081a081a00000000094c094c094c094c094c00000000004200420042000000000000000000000044f00000000000002100210021000000000000000160016001600000000000000004013000000000000000088118811881100000000000098009800000000000000000000004c1e00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004c1f0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
`endif

`ifdef RGB24
    `ifdef W128
        // this is abcdefghij placed in middle of displays
        // 2048 + 16
        localparam [(8*((384*3) + 2))-1:0] myled_row_basic = 'h4c04490229022902ab0acb02ec028a0a4a02280aa701a601a701a601a701c7010902ab128b0a0f4c9675346d9354d34c112c2d238b0a290a4a0a290a0902aa12ab12280aa7014501860186014501650186018609460145014501450125012401250124012501450145014501250145014501450125014501660186096601650166016501660186096601650946016501450144012501240125012401250124012501450125010401e4000301e400c3004601e300250144092501a611c711e719c811c719a7114a5b539d739d02090401e400e300a300a2008200820082008200620061006200610062006100620061006200810062008200820082008200a20083006501660186096601650946016501450144012501240125012401250124012501450125010401e4000301e400c3004601e300250144092501a611c711e719c811c719a7114a5b539d739d02090401e400e300a300a2008200820082008200620061006200610062006100620061006200810062008200820082008200a2008300490229022902ab0acb02ec028a0a4a02280aa701a601a701a601a701c7010902ab128b0a0f4c9675346d9354d34c112c2d238b0a290a4a0a290a0902aa12ab12280aa7014501860186014501650186018609460145014501450125012401250124012501450145014501250145014501450125014501660186096601650166016501660186096601650946016501450144012501240125012401250124012501450125010401e4000301e400c3004601e300250144092501a611c711e719c811c719a7114a5b539d739d02090401e400e300a300a2008200820082008200620061006200610062006100620061006200810062008200820082008200a20083006501660186096601650946016501450144012501240125012401250124012501450125010401e4000301e400c3004601e300250144092501a611c711e719c811c719a7114a5b539d739d02090401e400e300a300a2008200820082008200620061006200610062006100620061006200810062008200820082008200a2008300490229022902ab0acb02ec028a0a4a02280aa701a601a701a601a701c7010902ab128b0a0f4c9675346d9354d34c112c2d238b0a290a4a0a290a0902aa12ab12280aa7014501860186014501650186018609460145014501450125012401250124012501450145014501250145014501450125014501660186096601650166016501660186096601650946016501450144012501240125012401250124012501450125010401e4000301e400c3004601e300250144092501a611c711e719c811c719a7114a5b539d739d02090401e400e300a300a2008200820082008200620061006200610062006100620061006200810062008200820082008200a20083006501660186096601650946016501450144012501240125012401250124012501450125010401e4000301e400c3004601e300250144092501a611c711e719c811c719a7114a5b539d739d02090401e400e300a300a2008200820082008200620061006200610062006100620061006200810062008200820082008200a2008300;


    `else
        // 260 * 8 = 2080 ;; 64 * 2 * 8
        // 128 bytes (64 pixels * 2) * 8 bits + (1bytes * 8bits [L]) + (1bytes * 8bits [row]) == (64*2*8) + 8 + 8 = 1040
        // i don't know how we got to 260... pretty sure it should be 258.
        // 1024 + 16
        localparam [(8*((64*3) + 2))-1:0] myled_row_basic = 'h4c04_FFFEFD000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000_EFEEED;
        // FF-> 0x04fd (12bits)
        // FE-> 0x04fe
        // FD-> 0x04ff
        // EF-> 0x0401
        // EE-> 0x0402
        // ED-> 0x0403
    `endif
`else
    `ifdef W128
        // (2*256) + 2 = 514 * 8 = 4112
        // this is abcdefghij duplicated
        // logic [4111:0] myled_row = 'h4c040000000098000000000000009800000081a000000000000081a0000094c000000000000094c00000042000000000000004200000044f00000000000000000000021000000000000000000000001600000000000000160000401300000000000040130000000000008811000000000000000000000000980000000000000000000000000098000000000000009800000081a000000000000081a0000094c000000000000094c00000042000000000000004200000044f0000000000000000000002100000000000000000000000160000000000000016000040130000000000004013000000000000881100000000000000000000000098000000000000000000;
        // this is abcdefghij placed in middle of displays
        // 2048 + 16
        //              (PIXEL_WIDTH * COLOR_DEPTH) + (COMMAND + ROW)
        localparam [(8*((384*2) + 2))-1:0] myled_row_basic = 'h4c04490229022902ab0acb02ec028a0a4a02280aa701a601a701a601a701c7010902ab128b0a0f4c9675346d9354d34c112c2d238b0a290a4a0a290a0902aa12ab12280aa7014501860186014501650186018609460145014501450125012401250124012501450145014501250145014501450125014501660186096601650166016501660186096601650946016501450144012501240125012401250124012501450125010401e4000301e400c3004601e300250144092501a611c711e719c811c719a7114a5b539d739d02090401e400e300a300a2008200820082008200620061006200610062006100620061006200810062008200820082008200a2008300490229022902ab0acb02ec028a0a4a02280aa701a601a701a601a701c7010902ab128b0a0f4c9675346d9354d34c112c2d238b0a290a4a0a290a0902aa12ab12280aa701450186018601450165018601860946014501450145012501240125012401250145014501450125014501450145012501450166018609660165016601490229022902ab0acb02ec028a0a4a02280aa701a601a701a601a701c7010902ab128b0a0f4c9675346d9354d34c112c2d238b0a290a4a0a290a0902aa12ab12280aa7014501860186014501650186018609460145014501450125012401250124012501450145014501250145014501450125014501660186096601650166016501660186096601650946016501450144012501240125012401250124012501450125010401e4000301e400c3004601e300250144092501a611c711e719c811c719a7114a5b539d739d02090401e400e300a300a2008200820082008200620061006200610062006100620061006200810062008200820082008200a2008300490229022902ab0acb02ec028a0a4a02280aa701a601a701a601a701c7010902ab128b0a0f4c9675346d9354d34c112c2d238b0a290a4a0a290a0902aa12ab12280aa701450186018601450165018601860946014501450145012501240125012401250145014501450125014501450145012501450166018609660165016601;


    `else
        // 260 * 8 = 2080 ;; 64 * 2 * 8
        // 128 bytes (64 pixels * 2) * 8 bits + (1bytes * 8bits [L]) + (1bytes * 8bits [row]) == (64*2*8) + 8 + 8 = 1040
        // i don't know how we got to 260... pretty sure it should be 258.
        // 1024 + 16
        localparam [(8*((64*2) + 2))-1:0] myled_row_basic = 'h4c0449026b02cb0a6a02e7018701c701e801aa12d354345d5144cc1a4a02290a8b12c7016601850166016501450124012501440145014501450145014601650966016509660165014501440125012401250144010401e300040104014501c711c811a51971746c53a200c30082008200820061006200610062008200820082008300;
    `endif
`endif
// Add tests for pixel set command
localparam [(8*1)-1:0] myled_row_brightness_1 = 'h33; // "3"

localparam [(8*2)-1:0] myled_row_brightness_2 = 'h5423; // "T" + \x23
localparam [(8*2)-1:0] myled_row_brightness_3 = 'h5438; // "T" + \x38

localparam [(8*1)-1:0] myled_row_blankpanel = 'h5a;

`ifdef USE_WATCHDOG
    localparam [(8*(8+1))-1:0] myled_row_watchdog = 'h57_de_ad_be_ef_fe_eb_da_ed; // "W" + "DEADBEEFFEEBDAED"
`endif
`ifdef RGB24
    `ifdef W128
        localparam [(8*7)-1:0] myled_row_pixel  = 'h50_00_0078_132040; // "P" + row=8 column=0x30 bytedata=0x1020
        localparam [(8*7)-1:0] myled_row_pixel2 = 'h50_01_0079_304013;
        localparam [(8*4)-1:0] myled_row_fillpanel = 'h46_314287;
        localparam [(8*10)-1:0] myled_row_fillrect = 'h66_0001_0A_0071_05_E0A932; // "f" + x1/y1/width/height/color
    `else
        localparam [(8*6)-1:0] myled_row_pixel  = 'h50_00_30_132040; // "P" + row=8 column=0x30 bytedata=0x1020
        localparam [(8*6)-1:0] myled_row_pixel2 = 'h50_01_32_304013;
        localparam [(8*4)-1:0] myled_row_fillpanel = 'h46_314287;
        localparam [(8*8)-1:0] myled_row_fillrect = 'h66_05_0A_10_05_E0A932; // "f" + x1/y1/width/height/color
    `endif
`else
    `ifdef W128
        localparam [(8*6)-1:0] myled_row_pixel  = 'h50_00_0078_1020; // "P" + row=8 column=0x30 bytedata=0x1020
        localparam [(8*6)-1:0] myled_row_pixel2 = 'h50_01_0079_3040;
        localparam [(8*3)-1:0] myled_row_fillpanel = 'h46_3142;
        localparam [(8*9)-1:0] myled_row_fillrect = 'h66_0001_0A_0071_05_E0A9; // "f" + x1/y1/width/height/color
    `else
        localparam [(8*5)-1:0] myled_row_pixel  = 'h50_00_30_1020; // "P" + row=8 column=0x30 bytedata=0x1020
        localparam [(8*5)-1:0] myled_row_pixel2 = 'h50_01_32_3040;
        localparam [(8*3)-1:0] myled_row_fillpanel = 'h46_3142;
        localparam [(8*7)-1:0] myled_row_fillrect = 'h66_05_0A_10_05_E0A9; // "f" + x1/y1/width/height/color
    `endif
`endif
logic [
        ($bits(myled_row_blankpanel)
            + $bits(myled_row_fillpanel)
            + $bits(myled_row_fillrect)
            `ifdef USE_WATCHDOG
                + $bits(myled_row_watchdog)
            `endif
            `ifdef RGB24
                + $bits(myled_row_basic)
            `endif
            + $bits(myled_row_pixel)
            + $bits(myled_row_pixel2)
            + $bits(myled_row_brightness_1)
            + $bits(myled_row_brightness_2)
            + $bits(myled_row_brightness_3)
        )-1:0] myled_row = {
                                            myled_row_blankpanel,
                                            `ifdef USE_WATCHDOG
                                                myled_row_watchdog,
                                            `endif
                                            myled_row_fillpanel,
                                            myled_row_fillrect,
                                            myled_row_pixel,
                                            myled_row_pixel2,
                                            myled_row_brightness_1,
                                            myled_row_brightness_2,
                                            myled_row_brightness_3,
                                            myled_row_basic
                                        };

`ifdef JUNK
    //>>> "".join([a[i] for i in range(len(a)-1, -1, -1)])
    //'brR L-77665544332211887766554433221188776655443322118877665544332211887766554433221188776655443322118877665544332211887766554433221110'
    //logic [1071:0] mystring = "brR L-77665544332211887766554433221188776655443322118877665544332211887766554433221188776655443322118877665544332211887766554433221110";
    //logic [1071:0] mystring = 'h627252204c2d3737363635353434333332323131383837373636353534343333323231313838373736363535343433333232313138383737363635353434333332323131383837373636353534343333323231313838373736363535343433333232313138383737363635353434333332323131383837373636353534343333323231313130;
    //logic [2111:0] mystring = 'h627252204c2d37373636353534343333323231313838373736363535343433333232313138383737363635353434333332323131383837373636353534343333323231313838373736363535343433333232313138383737363635353434333332323131383837373636353534343333323231313838373736363535343433333232313131304c133737363635353434333332323131383837373636353534343333323231313838373736363535343433333232313138383737363635353434333332323131383837373636353534343333323231313838373736363535343433333232313138383737363635353434333332323131383837373636353534343333323231313130;

    // switched 4c18 to 4c09 (in an effort to align 4c09 with 4c19 [which immediately follows])
    // for some reason this seems to start simulating at 4c18 (row 22..)
    // also, for 4c09 added 0x1234 as first few pixels, and for 4c19 added 0x5678 for first few pixels
    // 8320 * 8 = 66560, log2=16.001... -> 17
    // mystring represents many concatenated led pixel rows (L01DATA,L02DATA...)
    // logic [66559:0] mystringfull = 'h4c0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004c0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004c0200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004c030000000000009800980098000000000081a081a081a081a000000000000094c094c094c000000000042004200420042000000000044f044f044f044f044f0000021002100210021002100000000000160016001600000000401300000000000040130000881188118811881188110000000000009800980098000000000000004c040000000098000000000000009800000081a000000000000081a0000094c000000000000094c00000042000000000000004200000044f00000000000000000000021000000000000000000000001600000000000000160000401300000000000040130000000000008811000000000000000000000000980000000000000000004c050000000098000000000000009800000081a000000000000081a0000094c000000000000000000000042000000000000004200000044f00000000000000000000021000000000000000000000001600000000000000000000401300000000000040130000000000008811000000000000000000000000980000000000000000004c060000000098000000000000009800000081a081a081a081a00000000094c000000000000000000000042000000000000004200000044f044f044f044f00000000021002100210021000000000001600000000000000000000401340134013401340130000000000008811000000000000000000000000980000000000000000004c070000000098009800980098009800000081a000000000000081a0000094c000000000000000000000042000000000000004200000044f00000000000000000000021000000000000000000000001600000000001600160000401300000000000040130000000000008811000000000000000000000000980000000000000000004c080000000098000000000000009800000081a000000000000081a0000094c000000000000094c00000042000000000000004200000044f00000000000000000000021000000000000000000000001600000000000000160000401300000000000040130000000000008811000000000000980000000000980000000000000000004c090000000098000000000000009800000081a081a081a081a000000000000094c094c094c000000000042004200420042000000000044f044f044f044f044f0000021000000000000000000000000000160016001600000000401300000000000040130000881188118811881188110000000098009800000000000000000000004c0a00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004c0b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004c0c00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004c0d00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004c0e0000000000000000000000000000000081a000000000000000000000000000000000000000000000000000000000000004200000000000000000000000000000000000000210021000000000000000000000000000000000401300000000000000000000000000008811000000000000000000000000980000000000000000004c0f0000000000000000000000000000000081a000000000000000000000000000000000000000000000000000000000000004200000000000000000000000000000000002100000000002100000000000000000000000000000401300000000000000000000000000000000000000000000000000000000000000000000000000004c100000000000009800980098000000000081a0000081a081a000000000000094c094c094c0000000000000042004200000042000000000044f044f044f00000000000002100000000000000000000000160016001600160000401300004013401300000000000000008811000000000000000000009800980000000000000000004c110000000000000000000000009800000081a081a00000000081a0000094c000000000000000000000042000000000042004200000044f000000000000044f0000021002100210000000000000001600000000000000160000401340130000000040130000000088118811000000000000000000000000980000000000000000004c120000000000009800980098009800000081a000000000000081a0000094c000000000000000000000042000000000000004200000044f044f044f044f00000000000002100000000000000000000000160016001600160000401300000000000040130000000000008811000000000000000000000000980000000000000000004c130000000098000000000000009800000081a000000000000081a0000094c000000000000094c00000042000000000000004200000044f00000000000000000000000002100000000000000000000000000000000000160000401300000000000040130000000000008811000000000000980000000000980000000000000000004c140000000000009800980098000000000081a081a081a081a000000000000094c094c094c0000000000000042004200420042000000000044f044f044f00000000000002100000000000000000000000160016001600000000401300000000000040130000000088118811881100000000000098009800000000000000000000004c1500000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004c1600000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004c17000000000000980098009800000000000000000081a0000000000000000094c094c094c000000000042004200420042004200000000000000000044f00000000021002100210021002100000000000000016001600000000401340134013401340130000000088118811881100000000000098009800980000000000000000004c0912340000980000000000000098000000000081a081a000000000000094c000000000000094c0000000000000000004200000000000000000044f044f00000000021000000000000000000000000000160000000000000000401300000000000040130000881100000000000088110000980000000000000098000000000000004c19567800009800000000009800980000000000000081a0000000000000000000000000000094c00000000000000420000000000000000002100000044f00000000021002100210021000000000001600000000000000000000000000000000401300000000881100000000000088110000980000000000000098000000000000004c1a000000009800000098000000980000000000000081a000000000000000000000000094c000000000000000000000042000000000044f00000000044f00000000000000000000000002100000001600160016001600000000000000000000401300000000000088118811881100000000000098009800980098000000000000004c1b000000009800980000000000980000000000000081a00000000000000000000094c0000000000000000000000000000004200000044f044f044f044f044f0000000000000000000002100000001600000000000000160000000000004013000000000000881100000000000088110000000000000000000098000000000000004c1c000000009800000000000000980000000000000081a0000000000000000094c00000000000000000042000000000000004200000000000000000044f00000000021000000000000002100000001600000000000000160000000000004013000000000000881100000000000088110000000000000000980000000000000000004c1d00000000000098009800980000000000000081a081a081a00000000094c094c094c094c094c00000000004200420042000000000000000000000044f00000000000002100210021000000000000000160016001600000000000000004013000000000000000088118811881100000000000098009800000000000000000000004c1e00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004c1f0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
`endif

`ifdef W128
    // (2*256) + 2 = 514 * 8 = 4112
    // this is abcdefghij duplicated
    // logic [4111:0] myled_row = 'h4c040000000098000000000000009800000081a000000000000081a0000094c000000000000094c00000042000000000000004200000044f00000000000000000000021000000000000000000000001600000000000000160000401300000000000040130000000000008811000000000000000000000000980000000000000000000000000098000000000000009800000081a000000000000081a0000094c000000000000094c00000042000000000000004200000044f0000000000000000000002100000000000000000000000160000000000000016000040130000000000004013000000000000881100000000000000000000000098000000000000000000;
    // this is abcdefghij placed in middle of displays
    localparam myled_row_size_basic = 2048 + 16;
    // See row4 of uart/w128_f60.uart
    logic [myled_row_size_basic-1:0] myled_row_basic = 'h4c04490229022902ab0acb02ec028a0a4a02280aa701a601a701a601a701c7010902ab128b0a0f4c9675346d9354d34c112c2d238b0a290a4a0a290a0902aa12ab12280aa7014501860186014501650186018609460145014501450125012401250124012501450145014501250145014501450125014501660186096601650166016501660186096601650946016501450144012501240125012401250124012501450125010401e4000301e400c3004601e300250144092501a611c711e719c811c719a7114a5b539d739d02090401e400e300a300a2008200820082008200620061006200610062006100620061006200810062008200820082008200a2008300;


`else
    // 260 * 8 = 2080 ;; 64 * 2 * 8
    // 128 bytes (64 pixels * 2) * 8 bits + (1bytes * 8bits [L]) + (1bytes * 8bits [row]) == (64*2*8) + 8 + 8 = 1040
    // i don't know how we got to 260... pretty sure it should be 258.
    localparam myled_row_size_basic = 1024 + 16;
    // See row4 of uart/w64_f60.uart
    logic [myled_row_size_basic-1:0] myled_row_basic = 'h4c0449026b02cb0a6a02e7018701c701e801aa12d354345d5144cc1a4a02290a8b12c7016601850166016501450124012501440145014501450145014601650966016509660165014501440125012401250144010401e300040104014501c711c811a51971746c53a200c30082008200820061006200610062008200820082008300;
;
`endif

// Add tests for pixel set command
localparam myled_row_size_pixel = (1 + 1 + 1 + 2) * 8;
logic [myled_row_size_pixel-1:0] myled_row_pixel  = 'h50_08_30_10_20;
logic [myled_row_size_pixel-1:0] myled_row_pixel2 = 'h50_09_32_30_40;


localparam myled_row_size = myled_row_size_basic + myled_row_size_pixel + myled_row_size_pixel;
logic [myled_row_size-1:0] myled_row = {myled_row_basic, myled_row_pixel, myled_row_pixel2};

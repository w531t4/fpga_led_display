module framebuffer_fetch (
	input reset,
	input clk_in,

	input [5:0] column_address,
	input [3:0] row_address,

	input pixel_load_start,

	input [15:0] ram_data_in,
	output [10:0] ram_address,
	output ram_clk_enable,
	output ram_reset,

	output reg [15:0] rgb565_top,
	output reg [15:0] rgb565_bottom,
	output [3:0] pixel_load_counter2
);
	wire ram_clk_enable_real;
	assign ram_clk_enable = ram_clk_enable_real;
	/* grab data on falling edge of pixel clock */
	//wire pixel_load_running;
`ifdef USE_FM6126A
	wire pixel_load_counter;
	assign pixel_load_counter2[3:0] = { 3'b0, pixel_load_counter };
`else
	wire [1:0] pixel_load_counter;
	assign pixel_load_counter2[3:0] = { 2'b0, pixel_load_counter[1:0] };
`endif

	reg half_address;
	assign ram_address = { half_address, row_address[3:0], ~column_address[5:0] };

	assign ram_reset = reset;

	timeout #(
`ifdef USE_FM6126A
		.COUNTER_WIDTH(1)
`else
		.COUNTER_WIDTH(2)
`endif
	) timeout_pixel_load (
		.reset(reset),
		.clk_in(clk_in),
		.start(pixel_load_start),
`ifdef USE_FM6126A
		.value(1'd1),
`else
		.value(2'd3),
`endif
		.counter(pixel_load_counter),
		.running(ram_clk_enable_real)
	)  /* synthesis syn_noprune=1 */  ;

	always @(negedge clk_in, posedge reset) begin
		if (reset) begin
			half_address <= 1'b0;

			rgb565_top    <= 16'd0;
			rgb565_bottom <= 16'd0;
		end
		else begin
`ifdef USE_FM6126A
			if (pixel_load_counter == 'd1) begin
				rgb565_top <= ram_data_in;
				half_address <= 1'b0;
			end
			else if (pixel_load_counter == 'd0) begin
				rgb565_bottom <= ram_data_in;
				half_address <= 1'b1;
			end
`else
			if (pixel_load_counter == 'd3) begin
				half_address <= 1'b0;
			end
			else if (pixel_load_counter == 'd2) begin
				half_address <= 1'b1;
			end
			else if (pixel_load_counter == 'd1) begin
				rgb565_top <= ram_data_in;
			end
			else if (pixel_load_counter == 'd0) begin
				rgb565_bottom <= ram_data_in;
			end
`endif
/*

			// the RAM requires _two_ clock cycles to read...
			 //  but change the address every clock cycle, so long as we respect the two-cycle fetch //
			if (pixel_load_counter == 'd3) begin
				// setup the top-half address //
				half_address <= 1'b0;
			end
			else if (pixel_load_counter == 'd2) begin
				// setup the bottom-half address //
				half_address <= 1'b1;
			end
			else if (pixel_load_counter == 'd1) begin
				// latch the pixel's value //
				rgb565_top <= ram_data_in;
			end
			else if (pixel_load_counter == 'd0) begin
				// latch the pixel's value //
				rgb565_bottom <= ram_data_in;
			end

			else begin
			end
			*/
		end
	end
endmodule

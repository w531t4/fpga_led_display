// SPDX-FileCopyrightText: 2025 Aaron White <w531t4@gmail.com>
// SPDX-License-Identifier: MIT
`default_nettype none
module control_cmd_fillrect #(
    // verilator lint_off UNUSEDPARAM
    parameter integer unsigned _UNUSED = 0
    // verilator lint_on UNUSEDPARAM
) (
    input reset,
    input [7:0] data_in,
    input enable,
    input clk,
    input mem_clk,

    output types::fb_addr_t addr,
    output logic [7:0] data_out,
    output logic ram_write_enable,
    output logic ram_access_start,
    output logic ready_for_data,
    output logic done
);
    localparam integer unsigned _NUM_COLUMN_BYTES_NEEDED = calc::num_bytes_to_contain($bits(types::col_addr_t));
    localparam types::col_addr_field_byte_index_t LAST_COL_BYTE_INDEX = types::col_addr_field_byte_index_t'(_NUM_COLUMN_BYTES_NEEDED - 1);
    typedef enum {
        STATE_X1_CAPTURE,      // 0
        STATE_Y1_CAPTURE,      // 1
        STATE_WIDTH_CAPTURE,   // 2
        STATE_HEIGHT_CAPTURE,  // 3
        STATE_COLOR_CAPTURE,   // 4
        STATE_START,           // 5
        STATE_RUNNING,         // 6
        STATE_PREDONE,         // 7
        STATE_DONE             // 8
    } ctrl_fsm_t;
    ctrl_fsm_t state;
    logic local_reset;
    // verilator lint_off UNUSEDSIGNAL
    types::col_addr_field_t x1;
    // TODO: This probably isn't the right type
    types::col_addr_field_t width;
    // verilator lint_on UNUSEDSIGNAL
    types::col_addr_field_byte_index_t x1_byte_counter;
    types::col_addr_field_byte_index_t width_byte_counter;
    types::row_addr_t y1;
    types::row_addr_count_t height;
    logic subcmd_enable;
    wire cmd_blankpanel_done;
    types::color_field_t selected_color;
    types::color_index_t capturebytes_remaining;


    logic done_inside, done_level;
    ff_sync #(
        .INIT_STATE(1'b0)
    ) done_sync (
        .clk(clk),
        .signal(done_inside),
        .reset(reset),
        .sync_level(done_level),
        .sync_pulse(done)
    );
    function automatic types::color_index_t reset_capturebytes_remaining();
        reset_capturebytes_remaining = types::color_index_t'(params::BYTES_PER_PIXEL - 1);
    endfunction
    always @(posedge clk) begin
        if (reset) begin
            subcmd_enable <= 1'b0;
            state <= STATE_X1_CAPTURE;
            done_inside <= 1'b0;
            ready_for_data <= 1'b1;
            capturebytes_remaining <= reset_capturebytes_remaining();
            selected_color <= 'b0;
            x1_byte_counter <= 'b0;
            width_byte_counter <= 'b0;
            x1 <= 'b0;
            width <= 'b0;
            y1 <= 'b0;
            height <= 'b0;
            local_reset <= 1'b0;
        end else begin
            case (state)
                STATE_X1_CAPTURE: begin
                    // Big Endian
                    if (enable) begin
                        x1.bytes[LAST_COL_BYTE_INDEX - x1_byte_counter] <= data_in;
                        if (x1_byte_counter == LAST_COL_BYTE_INDEX) begin
                            state <= STATE_Y1_CAPTURE;
                        end else x1_byte_counter <= x1_byte_counter + 1;
                    end
                end
                STATE_Y1_CAPTURE: begin
                    if (enable) begin
                        y1 <= types::row_addr_t'(data_in);
                        state <= STATE_WIDTH_CAPTURE;
                    end
                end
                STATE_WIDTH_CAPTURE: begin
                    // Big Endian
                    if (enable) begin
                        width.bytes[LAST_COL_BYTE_INDEX - width_byte_counter] <= data_in;
                        if (width_byte_counter == LAST_COL_BYTE_INDEX) begin
                            state <= STATE_HEIGHT_CAPTURE;
                        end else width_byte_counter <= width_byte_counter + 1;
                    end
                end
                STATE_HEIGHT_CAPTURE: begin
                    if (enable) begin
                        height <= types::row_addr_count_t'(data_in);
                        state <= STATE_COLOR_CAPTURE;
                        // The following assignment of width is done to reduce the burden on clk_root.
                        // TODO: types::col_addr_field_t' is the wrong type here - it's a _count_t that doesn't exist yet
                        width <= types::col_addr_field_t'(calc::clamp_remaining_dimension(
                            types::uint_t'(x1), types::uint_t'(width), params::PIXEL_WIDTH
                        ));
                    end
                end
                STATE_COLOR_CAPTURE: begin
                    // Big Endian
                    if (enable) begin
                        selected_color.bytes[capturebytes_remaining] <= data_in;
                        if (capturebytes_remaining == 0) begin
                            state <= STATE_START;
                            ready_for_data <= 1'b0;
                            // The following assignment of height is done to reduce the burden on clk_root.
                            height <= types::row_addr_count_t'(calc::clamp_remaining_dimension(
                                types::uint_t'(y1), types::uint_t'(height), params::PIXEL_HEIGHT
                            ));

                        end else begin
                            capturebytes_remaining <= capturebytes_remaining - 'd1;
                        end
                    end
                end
                STATE_START: begin
                    subcmd_enable <= 1'b1;
                    state <= STATE_RUNNING;
                end
                STATE_RUNNING: begin
                    if (cmd_blankpanel_done) begin
                        state <= STATE_PREDONE;
                        local_reset <= 1'b1;
                        subcmd_enable <= 1'b0;
                    end
                end
                STATE_PREDONE: begin
                    done_inside <= 1'b1;
                    local_reset <= 1'b0;
                    state <= STATE_DONE;
                end
                STATE_DONE: begin
                    done_inside <= 1'b0;
                    ready_for_data <= 1'b1;
                    state <= STATE_X1_CAPTURE;
                    x1_byte_counter <= 'b0;
                    width_byte_counter <= 'b0;
                    capturebytes_remaining <= reset_capturebytes_remaining();
                    selected_color <= 'b0;
                    x1 <= 'b0;
                    width <= 'b0;
                    y1 <= 'b0;
                    height <= 'b0;
                end
                default state <= state;
            endcase
        end
    end

    control_subcmd_fillarea #(
        ._UNUSED('d0)
    ) subcmd_fillarea (
        .reset(reset || local_reset),
        .enable(subcmd_enable),
        .clk(mem_clk),
        .ack(done),
        .x1(types::col_addr_t'(x1)),
        .y1(y1),
        .width(types::col_addr_count_t'(width)),
        .height(types::row_addr_count_t'(height)),
        .color(selected_color),
        .row(addr.row),
        .column(addr.col),
        .pixel(addr.pixel),
        .data_out(data_out),
        .ram_write_enable(ram_write_enable),
        .ram_access_start(ram_access_start),
        .done(cmd_blankpanel_done)
    );
    wire _unused_ok = &{1'b0, done_level, 1'b0};
endmodule

    // verilator lint_off UNUSEDPARAM
    parameter _NUM_SUBPANELS = PIXEL_HEIGHT / PIXEL_HALFHEIGHT,
    parameter _NUM_SUBPANELSELECT_BITS = $clog2(_NUM_SUBPANELS),
    parameter _NUM_PIXELCOLORSELECT_BITS = $clog2(BYTES_PER_PIXEL),
    parameter _NUM_ADDRESS_B_BITS = $clog2(PIXEL_HALFHEIGHT) + $clog2(PIXEL_WIDTH),
    parameter _NUM_ADDRESS_A_BITS = _NUM_SUBPANELSELECT_BITS + _NUM_PIXELCOLORSELECT_BITS + _NUM_ADDRESS_B_BITS,
    parameter _NUM_STRUCTURE_BITS = _NUM_ADDRESS_A_BITS - _NUM_ADDRESS_B_BITS,
    parameter _NUM_DATA_A_BITS = 8,
    parameter _NUM_DATA_B_BITS = ((1 << _NUM_PIXELCOLORSELECT_BITS) << _NUM_SUBPANELSELECT_BITS) << $clog2(8),
    parameter _NUM_BITS_PER_SUBPANEL = _NUM_DATA_B_BITS >> _NUM_SUBPANELSELECT_BITS,
    // verilator lint_on UNUSEDPARAM

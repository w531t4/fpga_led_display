parameter PIXEL_WIDTH = 64,
parameter PIXEL_HEIGHT = 32,
parameter PIXEL_HALFHEIGHT = 16,
parameter BYTES_PER_PIXEL = 2,

// SPDX-FileCopyrightText: 2025 Aaron White <w531t4@gmail.com>
// SPDX-License-Identifier: MIT
package types_pkg;
    typedef int unsigned uint_t;
endpackage

`timescale 1ns/100ps
module tb_main;
// context: RX DATA baud
// 16000000hz / 244444hz = 65.4547 ticks width=7
// tgt_hz variation (after rounding): 0.70%
// 16000000hz / 246154hz = 65 ticks width=7
parameter CTRLR_CLK_TICKS_PER_BIT = 7'd65;
parameter CTRLR_CLK_TICKS_WIDTH = 3'd7;


// context: TX DEBUG baud
// 16000000hz / 115200hz = 138.8889 ticks width=8
// tgt_hz variation (after rounding): -0.08%
// 16000000hz / 115108hz = 139 ticks width=8
parameter DEBUG_TX_UART_TICKS_PER_BIT = 8'd139;
parameter DEBUG_TX_UART_TICKS_PER_BIT_WIDTH = 4'd8;


// context: Debug msg rate
// 16000000hz / 22hz = 727272.7273 ticks width=20
// tgt_hz variation (after rounding): -0.00%
// 16000000hz / 22hz = 727273 ticks width=20
parameter DEBUG_MSGS_PER_SEC_TICKS = 20'd727273;
parameter DEBUG_MSGS_PER_SEC_TICKS_WIDTH = 5'd20;


`ifdef SIM
// use smaller value in testbench so we don't infinitely sim
parameter DEBUG_MSGS_PER_SEC_TICKS_SIM = 4'd15;
parameter DEBUG_MSGS_PER_SEC_TICKS_WIDTH_SIM = 3'd4;


// period = (1 / 16000000hz) / 2 = 31.25000
parameter SIM_HALF_PERIOD_NS = 31.25000;
`endif
    reg clk;
    wire clk_pixel;
    wire row_latch;
    wire OE;
    wire ROA0;
    wire ROA1;
    wire ROA2;
    wire ROA3;
    wire uart_rx;
    wire rgb2_0;
    wire rgb2_1;
    wire rbg2_2;
    wire rgb1_0;
    wire rgb1_1;
    wire rgb1_2;
    wire debugger_txout;
    reg  debugger_rxin;

    reg reset;
    reg local_reset;

    // debugger stuff
    wire debug_command_busy;
    wire debug_command_pulse;
    wire [7:0] debug_command;

    //>>> "".join([a[i] for i in range(len(a)-1, -1, -1)])
    //'brR L-77665544332211887766554433221188776655443322118877665544332211887766554433221188776655443322118877665544332211887766554433221110'
    //reg [1071:0] mystring = "brR L-77665544332211887766554433221188776655443322118877665544332211887766554433221188776655443322118877665544332211887766554433221110";
    //reg [1071:0] mystring = 'h627252204c2d3737363635353434333332323131383837373636353534343333323231313838373736363535343433333232313138383737363635353434333332323131383837373636353534343333323231313838373736363535343433333232313138383737363635353434333332323131383837373636353534343333323231313130;
    //reg [2111:0] mystring = 'h627252204c2d37373636353534343333323231313838373736363535343433333232313138383737363635353434333332323131383837373636353534343333323231313838373736363535343433333232313138383737363635353434333332323131383837373636353534343333323231313838373736363535343433333232313131304c133737363635353434333332323131383837373636353534343333323231313838373736363535343433333232313138383737363635353434333332323131383837373636353534343333323231313838373736363535343433333232313138383737363635353434333332323131383837373636353534343333323231313130;
    reg [8319:0] mystring = 'h4c0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004c0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004c0200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004c030000000000009800980098000000000081a081a081a081a000000000000094c094c094c000000000042004200420042000000000044f044f044f044f044f0000021002100210021002100000000000160016001600000000401300000000000040130000881188118811881188110000000000009800980098000000000000004c040000000098000000000000009800000081a000000000000081a0000094c000000000000094c00000042000000000000004200000044f00000000000000000000021000000000000000000000001600000000000000160000401300000000000040130000000000008811000000000000000000000000980000000000000000004c050000000098000000000000009800000081a000000000000081a0000094c000000000000000000000042000000000000004200000044f00000000000000000000021000000000000000000000001600000000000000000000401300000000000040130000000000008811000000000000000000000000980000000000000000004c060000000098000000000000009800000081a081a081a081a00000000094c000000000000000000000042000000000000004200000044f044f044f044f00000000021002100210021000000000001600000000000000000000401340134013401340130000000000008811000000000000000000000000980000000000000000004c070000000098009800980098009800000081a000000000000081a0000094c000000000000000000000042000000000000004200000044f00000000000000000000021000000000000000000000001600000000001600160000401300000000000040130000000000008811000000000000000000000000980000000000000000004c080000000098000000000000009800000081a000000000000081a0000094c000000000000094c00000042000000000000004200000044f00000000000000000000021000000000000000000000001600000000000000160000401300000000000040130000000000008811000000000000980000000000980000000000000000004c090000000098000000000000009800000081a081a081a081a000000000000094c094c094c000000000042004200420042000000000044f044f044f044f044f0000021000000000000000000000000000160016001600000000401300000000000040130000881188118811881188110000000098009800000000000000000000004c0a00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004c0b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004c0c00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004c0d00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004c0e0000000000000000000000000000000081a000000000000000000000000000000000000000000000000000000000000004200000000000000000000000000000000000000210021000000000000000000000000000000000401300000000000000000000000000008811000000000000000000000000980000000000000000004c0f0000000000000000000000000000000081a000000000000000000000000000000000000000000000000000000000000004200000000000000000000000000000000002100000000002100000000000000000000000000000401300000000000000000000000000000000000000000000000000000000000000000000000000004c100000000000009800980098000000000081a0000081a081a000000000000094c094c094c0000000000000042004200000042000000000044f044f044f00000000000002100000000000000000000000160016001600160000401300004013401300000000000000008811000000000000000000009800980000000000000000004c110000000000000000000000009800000081a081a00000000081a0000094c000000000000000000000042000000000042004200000044f000000000000044f0000021002100210000000000000001600000000000000160000401340130000000040130000000088118811000000000000000000000000980000000000000000004c120000000000009800980098009800000081a000000000000081a0000094c000000000000000000000042000000000000004200000044f044f044f044f00000000000002100000000000000000000000160016001600160000401300000000000040130000000000008811000000000000000000000000980000000000000000004c130000000098000000000000009800000081a000000000000081a0000094c000000000000094c00000042000000000000004200000044f00000000000000000000000002100000000000000000000000000000000000160000401300000000000040130000000000008811000000000000980000000000980000000000000000004c140000000000009800980098000000000081a081a081a081a000000000000094c094c094c0000000000000042004200420042000000000044f044f044f00000000000002100000000000000000000000160016001600000000401300000000000040130000000088118811881100000000000098009800000000000000000000004c1500000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004c1600000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004c17000000000000980098009800000000000000000081a0000000000000000094c094c094c000000000042004200420042004200000000000000000044f00000000021002100210021002100000000000000016001600000000401340134013401340130000000088118811881100000000000098009800980000000000000000004c1800000000980000000000000098000000000081a081a000000000000094c000000000000094c0000000000000000004200000000000000000044f044f00000000021000000000000000000000000000160000000000000000401300000000000040130000881100000000000088110000980000000000000098000000000000004c19000000009800000000009800980000000000000081a0000000000000000000000000000094c00000000000000420000000000000000002100000044f00000000021002100210021000000000001600000000000000000000000000000000401300000000881100000000000088110000980000000000000098000000000000004c1a000000009800000098000000980000000000000081a000000000000000000000000094c000000000000000000000042000000000044f00000000044f00000000000000000000000002100000001600160016001600000000000000000000401300000000000088118811881100000000000098009800980098000000000000004c1b000000009800980000000000980000000000000081a00000000000000000000094c0000000000000000000000000000004200000044f044f044f044f044f0000000000000000000002100000001600000000000000160000000000004013000000000000881100000000000088110000000000000000000098000000000000004c1c000000009800000000000000980000000000000081a0000000000000000094c00000000000000000042000000000000004200000000000000000044f00000000021000000000000002100000001600000000000000160000000000004013000000000000881100000000000088110000000000000000980000000000000000004c1d00000000000098009800980000000000000081a081a081a00000000094c094c094c094c094c00000000004200420042000000000000000000000044f00000000000002100210021000000000000000160016001600000000000000004013000000000000000088118811881100000000000098009800000000000000000000004c1e00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004c1f0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

    main tbi_main (
        .pin1(clk_pixel),
        .pin2(row_latch),
        .pin3(OE),
        .pin3_clk_16mhz(clk),
        .pin4(ROA0),
        .pin5(ROA1),
        .pin6(ROA2),
        .pin7(ROA3),
        .pin8(rgb1_0),
        .pin9(rgb1_1),
        .pin10(rgb1_2),
        .pin13(rgb2_2),
        .pin19(rgb2_0),
        .pin20(rgb2_1),
        .pin22(uart_rx),
        .pin23(debugger_txout),
        .pin24(debugger_rxin)
    );
    reg mask;
    debugger #(
		.DATA_WIDTH_BASE2(4'd14),
		.DATA_WIDTH(14'd8320),

        // use smaller than normal so it doesn't require us to simulate to
        // infinity to see results
		.DIVIDER_TICKS_WIDTH(DEBUG_MSGS_PER_SEC_TICKS_WIDTH_SIM),
		.DIVIDER_TICKS(DEBUG_MSGS_PER_SEC_TICKS_SIM),

		// We're using the debugger here as a data transmitter only. Need
		// to transmit at the same speed as the controller is expecting to
		// receive at
        .UART_TICKS_PER_BIT(CTRLR_CLK_TICKS_PER_BIT),
        .UART_TICKS_PER_BIT_SIZE(CTRLR_CLK_TICKS_WIDTH)
	) mydebug (
        .clk_in(clk && mask),
		.reset(local_reset),
		.data_in(mystring),
		.debug_uart_rx_in(1'b0),
		.debug_command(debug_command),
		.debug_command_pulse(debug_command_pulse),
		.debug_command_busy(debug_command_busy),
		.tx_out(uart_rx)
	);

    initial begin
        $dumpfile(`DUMP_FILE_NAME);
        $dumpvars(0, tb_main);
        clk = 0;
        mask = 0;


        debugger_rxin = 0;
        reset = 0;
        local_reset = 0;
        repeat (20) begin
            @(posedge clk);
        end
        @(posedge clk)
            local_reset = ! local_reset;
            reset = ! reset;
        @(posedge clk)
            local_reset = ! local_reset;
            reset = ! reset;
        repeat (20) begin
            @(posedge clk);
        end
        repeat (5) begin
            @(posedge clk);
        end
        @(posedge clk)
            mask = 1;
        #40000000 $finish;
    end
    always begin
        #SIM_HALF_PERIOD_NS clk <= !clk;
    end
endmodule

// SPDX-FileCopyrightText: 2025 Aaron White <w531t4@gmail.com>
// SPDX-License-Identifier: MIT
`ifndef SIM_DATA_SVH
`define SIM_DATA_SVH

// W384_RGB24_ROW_HEX:
//  - 9216 bits == 2304 characters == 1152 hex length
//  - 384 pixels (6x64)
`define W384_RGB24_ROW_HEX 'h490229022902ab0acb02ec028a0a4a02280aa701a601a701a601a701c7010902ab128b0a0f4c9675346d9354d34c112c2d238b0a290a4a0a290a0902aa12ab12280aa7014501860186014501650186018609460145014501450125012401250124012501450145014501250145014501450125014501660186096601650166016501660186096601650946016501450144012501240125012401250124012501450125010401e4000301e400c3004601e300250144092501a611c711e719c811c719a7114a5b539d739d02090401e400e300a300a2008200820082008200620061006200610062006100620061006200810062008200820082008200a20083006501660186096601650946016501450144012501240125012401250124012501450125010401e4000301e400c3004601e300250144092501a611c711e719c811c719a7114a5b539d739d02090401e400e300a300a2008200820082008200620061006200610062006100620061006200810062008200820082008200a2008300490229022902ab0acb02ec028a0a4a02280aa701a601a701a601a701c7010902ab128b0a0f4c9675346d9354d34c112c2d238b0a290a4a0a290a0902aa12ab12280aa7014501860186014501650186018609460145014501450125012401250124012501450145014501250145014501450125014501660186096601650166016501660186096601650946016501450144012501240125012401250124012501450125010401e4000301e400c3004601e300250144092501a611c711e719c811c719a7114a5b539d739d02090401e400e300a300a2008200820082008200620061006200610062006100620061006200810062008200820082008200a20083006501660186096601650946016501450144012501240125012401250124012501450125010401e4000301e400c3004601e300250144092501a611c711e719c811c719a7114a5b539d739d02090401e400e300a300a2008200820082008200620061006200610062006100620061006200810062008200820082008200a2008300490229022902ab0acb02ec028a0a4a02280aa701a601a701a601a701c7010902ab128b0a0f4c9675346d9354d34c112c2d238b0a290a4a0a290a0902aa12ab12280aa7014501860186014501650186018609460145014501450125012401250124012501450145014501250145014501450125014501660186096601650166016501660186096601650946016501450144012501240125012401250124012501450125010401e4000301e400c3004601e300250144092501a611c711e719c811c719a7114a5b539d739d02090401e400e300a300a2008200820082008200620061006200610062006100620061006200810062008200820082008200a20083006501660186096601650946016501450144012501240125012401250124012501450125010401e4000301e400c3004601e300250144092501a611c711e719c811c719a7114a5b539d739d02090401e400e300a300a2008200820082008200620061006200610062006100620061006200810062008200820082008200a2008300

// W64_RGB24_ROW_HEX:
//  - 1536 bits == 384 characters == 192 hex length
//  - 64 pixels (1x64)
`define W64_RGB24_ROW_HEX 'hFFFEFD000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000EFEEED
// FF-> 0x04fd (12bits)
// FE-> 0x04fe
// FD-> 0x04ff
// EF-> 0x0401
// EE-> 0x0402
// ED-> 0x0403

// W384_RGB565_ROW_HEX:
//  - 6144 bits == 1536 characters == 768 hex length
//  - 384 pixels (6x64)
`define W384_RGB565_ROW_HEX 'h490229022902ab0acb02ec028a0a4a02280aa701a601a701a601a701c7010902ab128b0a0f4c9675346d9354d34c112c2d238b0a290a4a0a290a0902aa12ab12280aa7014501860186014501650186018609460145014501450125012401250124012501450145014501250145014501450125014501660186096601650166016501660186096601650946016501450144012501240125012401250124012501450125010401e4000301e400c3004601e300250144092501a611c711e719c811c719a7114a5b539d739d02090401e400e300a300a2008200820082008200620061006200610062006100620061006200810062008200820082008200a2008300490229022902ab0acb02ec028a0a4a02280aa701a601a701a601a701c7010902ab128b0a0f4c9675346d9354d34c112c2d238b0a290a4a0a290a0902aa12ab12280aa701450186018601450165018601860946014501450145012501240125012401250145014501450125014501450145012501450166018609660165016601490229022902ab0acb02ec028a0a4a02280aa701a601a701a601a701c7010902ab128b0a0f4c9675346d9354d34c112c2d238b0a290a4a0a290a0902aa12ab12280aa7014501860186014501650186018609460145014501450125012401250124012501450145014501250145014501450125014501660186096601650166016501660186096601650946016501450144012501240125012401250124012501450125010401e4000301e400c3004601e300250144092501a611c711e719c811c719a7114a5b539d739d02090401e400e300a300a2008200820082008200620061006200610062006100620061006200810062008200820082008200a2008300490229022902ab0acb02ec028a0a4a02280aa701a601a701a601a701c7010902ab128b0a0f4c9675346d9354d34c112c2d238b0a290a4a0a290a0902aa12ab12280aa701450186018601450165018601860946014501450145012501240125012401250145014501450125014501450145012501450166018609660165016601

// W64_RGB565_ROW_HEX:
//  - 1024 bits == 256 characters == 128 hex length
//  - 64 pixels (1x64)
`define W64_RGB565_ROW_HEX 'h49026b02cb0a6a02e7018701c701e801aa12d354345d5144cc1a4a02290a8b12c7016601850166016501450124012501440145014501450145014601650966016509660165014501440125012401250144010401e300040104014501c711c811a51971746c53a200c30082008200820061006200610062008200820082008300

// Frame payload helpers: replicate the row sample across panel height.
// Cast to row_data_t so the row width (including leading zeros) is preserved.
`define W384_RGB24_FRAME_HEX  {params::PIXEL_HEIGHT{types::row_data_t'(`W384_RGB24_ROW_HEX)}}
`define W64_RGB24_FRAME_HEX   {params::PIXEL_HEIGHT{types::row_data_t'(`W64_RGB24_ROW_HEX)}}
`define W384_RGB565_FRAME_HEX {params::PIXEL_HEIGHT{types::row_data_t'(`W384_RGB565_ROW_HEX)}}
`define W64_RGB565_FRAME_HEX  {params::PIXEL_HEIGHT{types::row_data_t'(`W64_RGB565_ROW_HEX)}}

`endif

// SPDX-FileCopyrightText: 2025 Aaron White <w531t4@gmail.com>
// SPDX-License-Identifier: MIT
    // verilator lint_off UNUSEDPARAM
    localparam _NUM_SUBPANELS = PIXEL_HEIGHT / PIXEL_HALFHEIGHT,
    localparam _NUM_SUBPANELSELECT_BITS = $clog2(_NUM_SUBPANELS),
    localparam _NUM_PIXELCOLORSELECT_BITS = $clog2(params_pkg::BYTES_PER_PIXEL),
    localparam _NUM_COLUMN_ADDRESS_BITS = $clog2(PIXEL_WIDTH),
    localparam _NUM_ROW_ADDRESS_BITS = $clog2(PIXEL_HEIGHT),
    localparam _NUM_ADDRESS_B_BITS = $clog2(PIXEL_HALFHEIGHT) + _NUM_COLUMN_ADDRESS_BITS,
    localparam _NUM_ADDRESS_A_BITS = _NUM_SUBPANELSELECT_BITS + _NUM_PIXELCOLORSELECT_BITS + _NUM_ADDRESS_B_BITS,
    localparam _NUM_STRUCTURE_BITS = _NUM_ADDRESS_A_BITS - _NUM_ADDRESS_B_BITS,
    localparam _NUM_DATA_A_BITS = 8,
    localparam _NUM_DATA_B_BITS = ((1 << _NUM_PIXELCOLORSELECT_BITS) << _NUM_SUBPANELSELECT_BITS) << $clog2(8),
    localparam _NUM_BITS_PER_SUBPANEL = _NUM_DATA_B_BITS >> _NUM_SUBPANELSELECT_BITS,
    // verilator lint_on UNUSEDPARAM
